module tb_sfifo();
